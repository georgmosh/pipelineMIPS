library verilog;
use verilog.vl_types.all;
entity MyCircuit_vlg_vec_tst is
end MyCircuit_vlg_vec_tst;
