--REG_MEMWB.vhd
--This package implements a 16-bit pipeline register; using the behavioral MEM-WB register.
--Single structural operations are being implemented exploiting the logic from basic_func3.vhd
--All of the implemented operations in this file are styled in structural architecture.
--Authors: Georgios M. Moschovis (p3150113@aueb.gr)
--         Dimitrios Vetsis (p3120019@aueb.gr)

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

PACKAGE REG_MEMWB is

COMPONENT reg_MEM_WB
	GENERIC (n : INTEGER := 16);
	PORT (Result: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
				regAddress: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				Clock: IN STD_LOGIC;
				writeData: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
				writeAddress: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
		END COMPONENT;
		
END PACKAGE REG_MEMWB;

--package body declarations
LIBRARY ieee;
USE ieee.std_logic_1164.all;
--package body
ENTITY reg_MEM_WB IS 
	GENERIC (n : INTEGER := 16);
	PORT (Result: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
				regAddress: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				Clock: IN STD_LOGIC;
				writeData: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
				writeAddress: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END reg_MEM_WB;

ARCHITECTURE StructuralArchUnit OF reg_MEM_WB IS
	COMPONENT PipelineRegisterNo4 is
		GENERIC(n: INTEGER := 16);
		PORT (clk: IN STD_LOGIC;
				regaddress: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				res: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
				regaddressout: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
				out2: OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0));
	END COMPONENT;
	
	BEGIN
		    	--Component instantiations statements
		U0: PipelineRegisterNo4 PORT MAP(Clock, regAddress, Result, writeAddress, writeData);
END StructuralArchUnit;